`include "debug.vh"

module debug_tb;
    logic clk, rst;
    logic tck, tms, tdi, tdo;

endmodule
