`include "debug.vh"
`timescale 10ns/1ns
module debug_tb;
    // Want the period of clk over the period of tck to not be an
    // integer. This will test the synchronizers.
    int tcktime = 52;

    // DTM Signals
    logic clk, rst;
    logic tck, tms, tdi, tdo;
    dmi_t dmi_req;
    dmi_rsp_t dmi_rsp;

    dtm dut(
        clk, rst,
        tck, tms, tdi, tdo,
        dmi_req,
        dmi_rsp
    );

    initial begin
        tck = 1'b1;
        clk = 1'b1;
        forever #10 clk = ~clk; 
    end

    // Set of tasks to automate communicating over JTAG.
    task write_instr(input logic [4:0] INST);
        logic [11:0] tms_seq;
        logic [11:0] tdi_seq;
        begin
            tms_seq = {4'b0110, 5'b0, 3'b110};
            // Reverse instruction so LSB is first
            tdi_seq = {5'b0, {<<{INST}}, 2'b0};

            // Clock should be idling high, TMS should be low keeping
            // us in the Run-test/Idle state and the input should not
            // be driven.
            tck = 1;
            tms = 0;
            tdi = 0;
            
            // SelectIR -> CaptureIR -> ShiftIR
            for (int i = 11; i >= 0; i--) begin
                #(tcktime) tck = ~tck; // low
                tms = tms_seq[i];
                tdi = tdi_seq[i];
                #(tcktime) tck = ~tck; // high
            end
        end   
    endtask // instr

    // JTAG_DR Class that generalizes the task of reading and writing
    // to the Test Data Regisers. 
    class JTAG_DR #(parameter WIDTH = 32);
        task read(output logic [WIDTH-1:0] result);
            logic [5 + WIDTH + 2 - 1:0] tms_seq = {5'b01000, {(WIDTH-1){1'b0}}, 1'b1, 2'b10};
            for (int i = 5 + WIDTH + 2 - 1; i >= 0; i--) begin
                #(tcktime) tck = ~tck; 
                tdi = 0;
                tms = tms_seq[i];
                if ((i < WIDTH + 2) && (i >= 2))
                  $display(WIDTH - i + 2-1);
                    result[WIDTH - i + 2-1] = tdo;
                #(tcktime) tck = ~tck;
            end
        endtask
    endclass
    
    
    // Want the period of clk over the period of tck to not be an
    // integer. This will test the synchronizers.
    initial begin
        JTAG_DR #(32) idcode = new;
        JTAG_DR #(32) dtmcs = new;
        JTAG_DR #(32 + 2 + 7) dmireg = new;

        logic [31:0] idcode_result;
        logic [31:0] dtmcs_result;
        logic [32+2+7-1:0] dmi_result;
        
        rst = 0;
        tms = 1;
        @(posedge clk) tms = 0; rst = 1;
        @(negedge clk) rst = 0;

        // Read IDCODE
        write_instr(5'b00001);
        // read_datareg(data);
        idcode.read(idcode_result);
        
        assert(idcode_result == 32'h1002AC05) $display("Received IDCODE");
        else $display("IDCODE was corrupted.");

        test($bits(idcode_result));
        
        $stop;
    end
    
endmodule
